    ����          Assembly-CSharp   Menu+Position   xyz        pC=
�?  �C