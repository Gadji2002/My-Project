    ����          Assembly-CSharp   Menu+Position   xyz        pC=
�?  �C    ����          Assembly-CSharp   Menu+Rotation   xyz      �T߾   �   �